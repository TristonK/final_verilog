module getsec(
    input clk,
	 output reg clk_ls
);

reg [24:0] countclk;

initial
begin
   countclk=0;
	clk_ls=0;
end

always @(posedge clk)
 if(countclk==1250000)  
 begin
   countclk <=0;
   clk_ls <= ~clk_ls;
  end
 else
   countclk <= countclk+1;
	
endmodule 